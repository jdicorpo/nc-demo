module alu_16bit (overflow,
    zero,
    a,
    alu_control,
    b,
    result);
 output overflow;
 output zero;
 input [15:0] a;
 input [3:0] alu_control;
 input [15:0] b;
 output [15:0] result;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;

 sky130_fd_sc_hd__inv_2 _249_ (.A(net27),
    .Y(_204_));
 sky130_fd_sc_hd__inv_2 _250_ (.A(net6),
    .Y(_205_));
 sky130_fd_sc_hd__inv_2 _251_ (.A(net22),
    .Y(_206_));
 sky130_fd_sc_hd__inv_2 _252_ (.A(net14),
    .Y(_207_));
 sky130_fd_sc_hd__inv_2 _253_ (.A(net17),
    .Y(_208_));
 sky130_fd_sc_hd__and2b_1 _254_ (.A_N(net23),
    .B(net3),
    .X(_209_));
 sky130_fd_sc_hd__nand2b_1 _255_ (.A_N(net3),
    .B(net23),
    .Y(_210_));
 sky130_fd_sc_hd__nand2b_4 _256_ (.A_N(_209_),
    .B(_210_),
    .Y(_211_));
 sky130_fd_sc_hd__and2_4 _257_ (.A(net2),
    .B(net22),
    .X(_212_));
 sky130_fd_sc_hd__or2_4 _258_ (.A(net2),
    .B(net22),
    .X(_213_));
 sky130_fd_sc_hd__and2b_2 _259_ (.A_N(_212_),
    .B(_213_),
    .X(_214_));
 sky130_fd_sc_hd__inv_2 _260_ (.A(_214_),
    .Y(_215_));
 sky130_fd_sc_hd__nor2_1 _261_ (.A(_211_),
    .B(_214_),
    .Y(_216_));
 sky130_fd_sc_hd__and2b_1 _262_ (.A_N(net36),
    .B(net16),
    .X(_217_));
 sky130_fd_sc_hd__nand2b_2 _263_ (.A_N(net16),
    .B(net36),
    .Y(_218_));
 sky130_fd_sc_hd__nand2b_2 _264_ (.A_N(_217_),
    .B(_218_),
    .Y(_219_));
 sky130_fd_sc_hd__and2_1 _265_ (.A(net15),
    .B(net35),
    .X(_220_));
 sky130_fd_sc_hd__or2_1 _266_ (.A(net15),
    .B(net35),
    .X(_221_));
 sky130_fd_sc_hd__nand2b_2 _267_ (.A_N(_220_),
    .B(_221_),
    .Y(_222_));
 sky130_fd_sc_hd__or4b_4 _268_ (.A(_211_),
    .B(_219_),
    .C(_214_),
    .D_N(_222_),
    .X(_223_));
 sky130_fd_sc_hd__inv_2 _269_ (.A(_223_),
    .Y(_224_));
 sky130_fd_sc_hd__nand2_1 _270_ (.A(net7),
    .B(net27),
    .Y(_225_));
 sky130_fd_sc_hd__or2_1 _271_ (.A(net7),
    .B(net27),
    .X(_226_));
 sky130_fd_sc_hd__and2_1 _272_ (.A(_225_),
    .B(_226_),
    .X(_227_));
 sky130_fd_sc_hd__nand2_1 _273_ (.A(_225_),
    .B(_226_),
    .Y(_228_));
 sky130_fd_sc_hd__and2b_1 _274_ (.A_N(net25),
    .B(net5),
    .X(_229_));
 sky130_fd_sc_hd__nand2b_1 _275_ (.A_N(net25),
    .B(net5),
    .Y(_230_));
 sky130_fd_sc_hd__and2b_1 _276_ (.A_N(net5),
    .B(net25),
    .X(_231_));
 sky130_fd_sc_hd__nor2_1 _277_ (.A(_229_),
    .B(_231_),
    .Y(_232_));
 sky130_fd_sc_hd__nand2_1 _278_ (.A(net4),
    .B(net24),
    .Y(_233_));
 sky130_fd_sc_hd__or2_1 _279_ (.A(net4),
    .B(net24),
    .X(_234_));
 sky130_fd_sc_hd__nand2_2 _280_ (.A(_233_),
    .B(_234_),
    .Y(_235_));
 sky130_fd_sc_hd__or2_1 _281_ (.A(_205_),
    .B(net26),
    .X(_236_));
 sky130_fd_sc_hd__nand2_2 _282_ (.A(net6),
    .B(net26),
    .Y(_237_));
 sky130_fd_sc_hd__or2_1 _283_ (.A(net6),
    .B(net26),
    .X(_238_));
 sky130_fd_sc_hd__nand2_2 _284_ (.A(_237_),
    .B(_238_),
    .Y(_239_));
 sky130_fd_sc_hd__inv_2 _285_ (.A(_239_),
    .Y(_240_));
 sky130_fd_sc_hd__nand4_1 _286_ (.A(_228_),
    .B(_232_),
    .C(_235_),
    .D(_239_),
    .Y(_241_));
 sky130_fd_sc_hd__or2_4 _287_ (.A(_223_),
    .B(_241_),
    .X(_242_));
 sky130_fd_sc_hd__and2_1 _288_ (.A(net12),
    .B(net32),
    .X(_243_));
 sky130_fd_sc_hd__xor2_4 _289_ (.A(net12),
    .B(net32),
    .X(_244_));
 sky130_fd_sc_hd__xnor2_1 _290_ (.A(net12),
    .B(net32),
    .Y(_245_));
 sky130_fd_sc_hd__or2_1 _291_ (.A(net13),
    .B(net33),
    .X(_246_));
 sky130_fd_sc_hd__nand2_1 _292_ (.A(net13),
    .B(net33),
    .Y(_247_));
 sky130_fd_sc_hd__xor2_2 _293_ (.A(net13),
    .B(net33),
    .X(_248_));
 sky130_fd_sc_hd__nand2_1 _294_ (.A(_246_),
    .B(_247_),
    .Y(_000_));
 sky130_fd_sc_hd__nor2_1 _295_ (.A(net11),
    .B(net31),
    .Y(_001_));
 sky130_fd_sc_hd__and2_1 _296_ (.A(net11),
    .B(net31),
    .X(_002_));
 sky130_fd_sc_hd__nor2_1 _297_ (.A(_001_),
    .B(_002_),
    .Y(_003_));
 sky130_fd_sc_hd__or2_1 _298_ (.A(net14),
    .B(net34),
    .X(_004_));
 sky130_fd_sc_hd__xor2_4 _299_ (.A(net14),
    .B(net34),
    .X(_005_));
 sky130_fd_sc_hd__nor2_1 _300_ (.A(_248_),
    .B(_005_),
    .Y(_006_));
 sky130_fd_sc_hd__or3b_4 _301_ (.A(_244_),
    .B(_003_),
    .C_N(_006_),
    .X(_007_));
 sky130_fd_sc_hd__and2b_1 _302_ (.A_N(net30),
    .B(net10),
    .X(_008_));
 sky130_fd_sc_hd__or2_1 _303_ (.A(net10),
    .B(net30),
    .X(_009_));
 sky130_fd_sc_hd__xnor2_2 _304_ (.A(net10),
    .B(net30),
    .Y(_010_));
 sky130_fd_sc_hd__and2b_1 _305_ (.A_N(net29),
    .B(net9),
    .X(_011_));
 sky130_fd_sc_hd__and2_4 _306_ (.A(net9),
    .B(net29),
    .X(_012_));
 sky130_fd_sc_hd__nor2_1 _307_ (.A(net9),
    .B(net29),
    .Y(_013_));
 sky130_fd_sc_hd__nor2_1 _308_ (.A(_012_),
    .B(_013_),
    .Y(_014_));
 sky130_fd_sc_hd__xnor2_1 _309_ (.A(net9),
    .B(net29),
    .Y(_015_));
 sky130_fd_sc_hd__and2_1 _310_ (.A(_010_),
    .B(_015_),
    .X(_016_));
 sky130_fd_sc_hd__and2b_1 _311_ (.A_N(net28),
    .B(net8),
    .X(_017_));
 sky130_fd_sc_hd__or2_1 _312_ (.A(net8),
    .B(net28),
    .X(_018_));
 sky130_fd_sc_hd__nand2_1 _313_ (.A(net8),
    .B(net28),
    .Y(_019_));
 sky130_fd_sc_hd__xnor2_4 _314_ (.A(net28),
    .B(net8),
    .Y(_020_));
 sky130_fd_sc_hd__nand2b_1 _315_ (.A_N(net1),
    .B(net21),
    .Y(_021_));
 sky130_fd_sc_hd__a21o_1 _316_ (.A1(_020_),
    .A2(_021_),
    .B1(_017_),
    .X(_022_));
 sky130_fd_sc_hd__nand2_1 _317_ (.A(_016_),
    .B(_022_),
    .Y(_023_));
 sky130_fd_sc_hd__a21o_1 _318_ (.A1(_010_),
    .A2(_011_),
    .B1(_008_),
    .X(_024_));
 sky130_fd_sc_hd__a21oi_2 _319_ (.A1(_016_),
    .A2(_022_),
    .B1(_024_),
    .Y(_025_));
 sky130_fd_sc_hd__and2b_1 _320_ (.A_N(net32),
    .B(net12),
    .X(_026_));
 sky130_fd_sc_hd__and2b_1 _321_ (.A_N(net31),
    .B(net11),
    .X(_027_));
 sky130_fd_sc_hd__a21o_1 _322_ (.A1(_245_),
    .A2(_027_),
    .B1(_026_),
    .X(_028_));
 sky130_fd_sc_hd__nand2b_1 _323_ (.A_N(net33),
    .B(net13),
    .Y(_029_));
 sky130_fd_sc_hd__or2_1 _324_ (.A(_005_),
    .B(_029_),
    .X(_030_));
 sky130_fd_sc_hd__o2bb2a_1 _325_ (.A1_N(_028_),
    .A2_N(_006_),
    .B1(net34),
    .B2(_207_),
    .X(_031_));
 sky130_fd_sc_hd__o211ai_4 _326_ (.A1(_007_),
    .A2(_025_),
    .B1(_030_),
    .C1(_031_),
    .Y(_032_));
 sky130_fd_sc_hd__nand2b_1 _327_ (.A_N(net15),
    .B(net35),
    .Y(_033_));
 sky130_fd_sc_hd__a21o_1 _328_ (.A1(_218_),
    .A2(_033_),
    .B1(_217_),
    .X(_034_));
 sky130_fd_sc_hd__o21a_1 _329_ (.A1(net2),
    .A2(_206_),
    .B1(_210_),
    .X(_035_));
 sky130_fd_sc_hd__o32a_1 _330_ (.A1(_211_),
    .A2(net57),
    .A3(_034_),
    .B1(_035_),
    .B2(_209_),
    .X(_036_));
 sky130_fd_sc_hd__and2b_1 _331_ (.A_N(net4),
    .B(net24),
    .X(_037_));
 sky130_fd_sc_hd__o211a_1 _332_ (.A1(_231_),
    .A2(_037_),
    .B1(_239_),
    .C1(_230_),
    .X(_038_));
 sky130_fd_sc_hd__a21oi_1 _333_ (.A1(_205_),
    .A2(net26),
    .B1(_038_),
    .Y(_039_));
 sky130_fd_sc_hd__o211a_1 _334_ (.A1(_241_),
    .A2(_036_),
    .B1(_039_),
    .C1(_228_),
    .X(_040_));
 sky130_fd_sc_hd__o21ai_1 _335_ (.A1(_242_),
    .A2(_032_),
    .B1(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__nand2_1 _336_ (.A(net1),
    .B(net21),
    .Y(_042_));
 sky130_fd_sc_hd__or2_1 _337_ (.A(net1),
    .B(net21),
    .X(_043_));
 sky130_fd_sc_hd__nand2_1 _338_ (.A(_042_),
    .B(_043_),
    .Y(_044_));
 sky130_fd_sc_hd__and3_1 _339_ (.A(_016_),
    .B(_020_),
    .C(_044_),
    .X(_045_));
 sky130_fd_sc_hd__or3b_1 _340_ (.A(_242_),
    .B(_007_),
    .C_N(_045_),
    .X(_046_));
 sky130_fd_sc_hd__nor2_1 _341_ (.A(net18),
    .B(net20),
    .Y(_047_));
 sky130_fd_sc_hd__o2111a_1 _342_ (.A1(net7),
    .A2(_204_),
    .B1(net17),
    .C1(net19),
    .D1(_047_),
    .X(_048_));
 sky130_fd_sc_hd__nor3b_1 _343_ (.A(net20),
    .B(net19),
    .C_N(net18),
    .Y(_049_));
 sky130_fd_sc_hd__or3b_4 _344_ (.A(net20),
    .B(net19),
    .C_N(net18),
    .X(_050_));
 sky130_fd_sc_hd__nand2_1 _345_ (.A(_208_),
    .B(_042_),
    .Y(_051_));
 sky130_fd_sc_hd__and3_2 _346_ (.A(_208_),
    .B(net19),
    .C(_047_),
    .X(_052_));
 sky130_fd_sc_hd__or4b_1 _347_ (.A(net17),
    .B(net18),
    .C(net20),
    .D_N(net19),
    .X(_053_));
 sky130_fd_sc_hd__or3_2 _348_ (.A(net18),
    .B(net20),
    .C(net19),
    .X(_054_));
 sky130_fd_sc_hd__a21oi_1 _349_ (.A1(net55),
    .A2(_054_),
    .B1(_044_),
    .Y(_055_));
 sky130_fd_sc_hd__a31o_1 _350_ (.A1(_041_),
    .A2(_046_),
    .A3(_048_),
    .B1(_055_),
    .X(_056_));
 sky130_fd_sc_hd__a31o_1 _351_ (.A1(_043_),
    .A2(net56),
    .A3(_051_),
    .B1(_056_),
    .X(net38));
 sky130_fd_sc_hd__nor2_4 _352_ (.A(_208_),
    .B(_050_),
    .Y(_057_));
 sky130_fd_sc_hd__nor2_4 _353_ (.A(net17),
    .B(_054_),
    .Y(_058_));
 sky130_fd_sc_hd__or2_2 _354_ (.A(net17),
    .B(_054_),
    .X(_059_));
 sky130_fd_sc_hd__or2_4 _355_ (.A(_020_),
    .B(_042_),
    .X(_060_));
 sky130_fd_sc_hd__nand2_1 _356_ (.A(_020_),
    .B(_042_),
    .Y(_061_));
 sky130_fd_sc_hd__nor2_2 _357_ (.A(_208_),
    .B(_054_),
    .Y(_062_));
 sky130_fd_sc_hd__or2_4 _358_ (.A(_208_),
    .B(_054_),
    .X(_063_));
 sky130_fd_sc_hd__a21oi_1 _359_ (.A1(_020_),
    .A2(_021_),
    .B1(_063_),
    .Y(_064_));
 sky130_fd_sc_hd__o21a_1 _360_ (.A1(_020_),
    .A2(_021_),
    .B1(_064_),
    .X(_065_));
 sky130_fd_sc_hd__o22a_1 _361_ (.A1(_019_),
    .A2(_050_),
    .B1(net55),
    .B2(_020_),
    .X(_066_));
 sky130_fd_sc_hd__a32o_1 _362_ (.A1(_058_),
    .A2(_060_),
    .A3(_061_),
    .B1(_057_),
    .B2(_018_),
    .X(_067_));
 sky130_fd_sc_hd__or3b_4 _363_ (.A(_067_),
    .B(_065_),
    .C_N(_066_),
    .X(net45));
 sky130_fd_sc_hd__o21ai_4 _364_ (.A1(_042_),
    .A2(_020_),
    .B1(_019_),
    .Y(_068_));
 sky130_fd_sc_hd__xnor2_1 _365_ (.A(_014_),
    .B(_068_),
    .Y(_069_));
 sky130_fd_sc_hd__nor2_1 _366_ (.A(_015_),
    .B(_022_),
    .Y(_070_));
 sky130_fd_sc_hd__a21o_1 _367_ (.A1(_015_),
    .A2(_022_),
    .B1(_063_),
    .X(_071_));
 sky130_fd_sc_hd__nor2_1 _368_ (.A(net17),
    .B(_012_),
    .Y(_072_));
 sky130_fd_sc_hd__o22a_1 _369_ (.A1(_012_),
    .A2(net55),
    .B1(_072_),
    .B2(_050_),
    .X(_073_));
 sky130_fd_sc_hd__o22a_1 _370_ (.A1(_059_),
    .A2(_069_),
    .B1(_070_),
    .B2(_071_),
    .X(_074_));
 sky130_fd_sc_hd__o21ai_1 _371_ (.A1(_013_),
    .A2(_073_),
    .B1(_074_),
    .Y(net46));
 sky130_fd_sc_hd__a21o_1 _372_ (.A1(_014_),
    .A2(_068_),
    .B1(_012_),
    .X(_075_));
 sky130_fd_sc_hd__xnor2_1 _373_ (.A(_010_),
    .B(_075_),
    .Y(_076_));
 sky130_fd_sc_hd__a211o_1 _374_ (.A1(_015_),
    .A2(_022_),
    .B1(_010_),
    .C1(_011_),
    .X(_077_));
 sky130_fd_sc_hd__a21oi_1 _375_ (.A1(_010_),
    .A2(_011_),
    .B1(_063_),
    .Y(_078_));
 sky130_fd_sc_hd__and3_1 _376_ (.A(_023_),
    .B(_077_),
    .C(_078_),
    .X(_079_));
 sky130_fd_sc_hd__nor2_1 _377_ (.A(_010_),
    .B(net55),
    .Y(_080_));
 sky130_fd_sc_hd__and3_1 _378_ (.A(net10),
    .B(net30),
    .C(net56),
    .X(_081_));
 sky130_fd_sc_hd__a211o_1 _379_ (.A1(_009_),
    .A2(_057_),
    .B1(_080_),
    .C1(_081_),
    .X(_082_));
 sky130_fd_sc_hd__a211o_1 _380_ (.A1(_058_),
    .A2(_076_),
    .B1(_082_),
    .C1(_079_),
    .X(net47));
 sky130_fd_sc_hd__a221o_1 _381_ (.A1(net10),
    .A2(net30),
    .B1(_068_),
    .B2(_014_),
    .C1(_012_),
    .X(_083_));
 sky130_fd_sc_hd__and3_1 _382_ (.A(_003_),
    .B(_083_),
    .C(_009_),
    .X(_084_));
 sky130_fd_sc_hd__a21oi_1 _383_ (.A1(_009_),
    .A2(_083_),
    .B1(_003_),
    .Y(_085_));
 sky130_fd_sc_hd__nor2_1 _384_ (.A(net17),
    .B(_002_),
    .Y(_086_));
 sky130_fd_sc_hd__o22a_1 _385_ (.A1(_002_),
    .A2(net55),
    .B1(_086_),
    .B2(_050_),
    .X(_087_));
 sky130_fd_sc_hd__and2_1 _386_ (.A(_003_),
    .B(_025_),
    .X(_088_));
 sky130_fd_sc_hd__nor2_1 _387_ (.A(_003_),
    .B(_025_),
    .Y(_089_));
 sky130_fd_sc_hd__o32a_1 _388_ (.A1(_063_),
    .A2(_088_),
    .A3(_089_),
    .B1(_087_),
    .B2(_001_),
    .X(_090_));
 sky130_fd_sc_hd__o31ai_1 _389_ (.A1(_059_),
    .A2(_084_),
    .A3(_085_),
    .B1(_090_),
    .Y(net48));
 sky130_fd_sc_hd__o21ai_1 _390_ (.A1(_027_),
    .A2(_089_),
    .B1(_245_),
    .Y(_091_));
 sky130_fd_sc_hd__nor3_1 _391_ (.A(_244_),
    .B(_003_),
    .C(_025_),
    .Y(_092_));
 sky130_fd_sc_hd__o311a_1 _392_ (.A1(_245_),
    .A2(_027_),
    .A3(_089_),
    .B1(_091_),
    .C1(_062_),
    .X(_093_));
 sky130_fd_sc_hd__o21a_1 _393_ (.A1(net12),
    .A2(net32),
    .B1(_057_),
    .X(_094_));
 sky130_fd_sc_hd__a221o_1 _394_ (.A1(_243_),
    .A2(net56),
    .B1(_052_),
    .B2(_244_),
    .C1(_094_),
    .X(_095_));
 sky130_fd_sc_hd__o21ai_1 _395_ (.A1(_002_),
    .A2(_084_),
    .B1(_244_),
    .Y(_096_));
 sky130_fd_sc_hd__o311a_1 _396_ (.A1(_244_),
    .A2(_002_),
    .A3(_084_),
    .B1(_096_),
    .C1(_058_),
    .X(_097_));
 sky130_fd_sc_hd__or3_4 _397_ (.A(_093_),
    .B(_095_),
    .C(_097_),
    .X(net49));
 sky130_fd_sc_hd__or3_1 _398_ (.A(_000_),
    .B(_028_),
    .C(_092_),
    .X(_098_));
 sky130_fd_sc_hd__o21ai_1 _399_ (.A1(_028_),
    .A2(_092_),
    .B1(_000_),
    .Y(_099_));
 sky130_fd_sc_hd__a21o_1 _400_ (.A1(_244_),
    .A2(_002_),
    .B1(_243_),
    .X(_100_));
 sky130_fd_sc_hd__a21oi_1 _401_ (.A1(_244_),
    .A2(_084_),
    .B1(_100_),
    .Y(_101_));
 sky130_fd_sc_hd__xnor2_1 _402_ (.A(_248_),
    .B(_101_),
    .Y(_102_));
 sky130_fd_sc_hd__nand2_1 _403_ (.A(_208_),
    .B(_247_),
    .Y(_103_));
 sky130_fd_sc_hd__a32o_1 _404_ (.A1(_246_),
    .A2(net56),
    .A3(_103_),
    .B1(_052_),
    .B2(_248_),
    .X(_104_));
 sky130_fd_sc_hd__a31o_1 _405_ (.A1(_062_),
    .A2(_098_),
    .A3(_099_),
    .B1(_104_),
    .X(_105_));
 sky130_fd_sc_hd__a21o_1 _406_ (.A1(_058_),
    .A2(_102_),
    .B1(_105_),
    .X(net50));
 sky130_fd_sc_hd__a21oi_1 _407_ (.A1(_029_),
    .A2(_099_),
    .B1(_005_),
    .Y(_106_));
 sky130_fd_sc_hd__a31o_1 _408_ (.A1(_005_),
    .A2(_029_),
    .A3(_099_),
    .B1(_063_),
    .X(_107_));
 sky130_fd_sc_hd__nor2_1 _409_ (.A(_106_),
    .B(_107_),
    .Y(_108_));
 sky130_fd_sc_hd__o21ai_1 _410_ (.A1(_000_),
    .A2(_101_),
    .B1(_247_),
    .Y(_109_));
 sky130_fd_sc_hd__xor2_1 _411_ (.A(_005_),
    .B(_109_),
    .X(_110_));
 sky130_fd_sc_hd__and3_1 _412_ (.A(net14),
    .B(net34),
    .C(net56),
    .X(_111_));
 sky130_fd_sc_hd__a221o_1 _413_ (.A1(_005_),
    .A2(_052_),
    .B1(_057_),
    .B2(_004_),
    .C1(_111_),
    .X(_112_));
 sky130_fd_sc_hd__a211o_1 _414_ (.A1(_058_),
    .A2(_110_),
    .B1(_112_),
    .C1(_108_),
    .X(net51));
 sky130_fd_sc_hd__and2_1 _415_ (.A(_248_),
    .B(_005_),
    .X(_113_));
 sky130_fd_sc_hd__and3_1 _416_ (.A(_244_),
    .B(_003_),
    .C(_113_),
    .X(_114_));
 sky130_fd_sc_hd__o211a_1 _417_ (.A1(net14),
    .A2(net34),
    .B1(net13),
    .C1(net33),
    .X(_115_));
 sky130_fd_sc_hd__a21oi_1 _418_ (.A1(net14),
    .A2(net34),
    .B1(_115_),
    .Y(_116_));
 sky130_fd_sc_hd__and2_1 _419_ (.A(_100_),
    .B(_113_),
    .X(_117_));
 sky130_fd_sc_hd__a31oi_2 _420_ (.A1(_009_),
    .A2(net58),
    .A3(_114_),
    .B1(_117_),
    .Y(_118_));
 sky130_fd_sc_hd__a21oi_2 _421_ (.A1(_116_),
    .A2(_118_),
    .B1(_222_),
    .Y(_119_));
 sky130_fd_sc_hd__a31o_1 _422_ (.A1(_222_),
    .A2(_116_),
    .A3(_118_),
    .B1(_059_),
    .X(_120_));
 sky130_fd_sc_hd__nor2_1 _423_ (.A(_222_),
    .B(_032_),
    .Y(_121_));
 sky130_fd_sc_hd__and2_1 _424_ (.A(_222_),
    .B(_032_),
    .X(_122_));
 sky130_fd_sc_hd__or3_1 _425_ (.A(_063_),
    .B(_121_),
    .C(_122_),
    .X(_123_));
 sky130_fd_sc_hd__o21ai_1 _426_ (.A1(net17),
    .A2(_220_),
    .B1(_221_),
    .Y(_124_));
 sky130_fd_sc_hd__o22a_1 _427_ (.A1(_222_),
    .A2(net55),
    .B1(_119_),
    .B2(_120_),
    .X(_125_));
 sky130_fd_sc_hd__o211ai_1 _428_ (.A1(_050_),
    .A2(_124_),
    .B1(_125_),
    .C1(_123_),
    .Y(net52));
 sky130_fd_sc_hd__o21ai_1 _429_ (.A1(_220_),
    .A2(_119_),
    .B1(_219_),
    .Y(_126_));
 sky130_fd_sc_hd__or3_1 _430_ (.A(_219_),
    .B(_220_),
    .C(_119_),
    .X(_127_));
 sky130_fd_sc_hd__and2b_1 _431_ (.A_N(net35),
    .B(net15),
    .X(_128_));
 sky130_fd_sc_hd__a21o_1 _432_ (.A1(_222_),
    .A2(_032_),
    .B1(_128_),
    .X(_129_));
 sky130_fd_sc_hd__xnor2_1 _433_ (.A(_219_),
    .B(_129_),
    .Y(_130_));
 sky130_fd_sc_hd__or2_1 _434_ (.A(net16),
    .B(net36),
    .X(_131_));
 sky130_fd_sc_hd__and2_1 _435_ (.A(net16),
    .B(net36),
    .X(_132_));
 sky130_fd_sc_hd__nand2_1 _436_ (.A(net16),
    .B(net36),
    .Y(_133_));
 sky130_fd_sc_hd__nor2_1 _437_ (.A(net55),
    .B(_132_),
    .Y(_134_));
 sky130_fd_sc_hd__o21a_1 _438_ (.A1(_057_),
    .A2(_134_),
    .B1(_131_),
    .X(_135_));
 sky130_fd_sc_hd__a221o_1 _439_ (.A1(_062_),
    .A2(_130_),
    .B1(_132_),
    .B2(net56),
    .C1(_135_),
    .X(_136_));
 sky130_fd_sc_hd__a31o_1 _440_ (.A1(_058_),
    .A2(_126_),
    .A3(_127_),
    .B1(_136_),
    .X(net53));
 sky130_fd_sc_hd__o31a_1 _441_ (.A1(_220_),
    .A2(_119_),
    .A3(_132_),
    .B1(_131_),
    .X(_137_));
 sky130_fd_sc_hd__xnor2_1 _442_ (.A(_215_),
    .B(_137_),
    .Y(_138_));
 sky130_fd_sc_hd__o31a_1 _443_ (.A1(net59),
    .A2(_122_),
    .A3(_128_),
    .B1(_218_),
    .X(_139_));
 sky130_fd_sc_hd__or2_1 _444_ (.A(_215_),
    .B(_139_),
    .X(_140_));
 sky130_fd_sc_hd__o311ai_2 _445_ (.A1(net59),
    .A2(_122_),
    .A3(_128_),
    .B1(_218_),
    .C1(_215_),
    .Y(_141_));
 sky130_fd_sc_hd__and3_1 _446_ (.A(_062_),
    .B(_140_),
    .C(_141_),
    .X(_142_));
 sky130_fd_sc_hd__o211a_1 _447_ (.A1(net17),
    .A2(_212_),
    .B1(_213_),
    .C1(net56),
    .X(_143_));
 sky130_fd_sc_hd__a22o_1 _448_ (.A1(_214_),
    .A2(_052_),
    .B1(_058_),
    .B2(_138_),
    .X(_144_));
 sky130_fd_sc_hd__or3_1 _449_ (.A(_142_),
    .B(_143_),
    .C(_144_),
    .X(net39));
 sky130_fd_sc_hd__a21oi_1 _450_ (.A1(_214_),
    .A2(_137_),
    .B1(_212_),
    .Y(_145_));
 sky130_fd_sc_hd__xnor2_1 _451_ (.A(_211_),
    .B(_145_),
    .Y(_146_));
 sky130_fd_sc_hd__nand2_1 _452_ (.A(net2),
    .B(_206_),
    .Y(_147_));
 sky130_fd_sc_hd__a21oi_1 _453_ (.A1(_141_),
    .A2(_147_),
    .B1(_211_),
    .Y(_148_));
 sky130_fd_sc_hd__a31o_1 _454_ (.A1(_211_),
    .A2(_141_),
    .A3(_147_),
    .B1(_063_),
    .X(_149_));
 sky130_fd_sc_hd__nor2_1 _455_ (.A(_148_),
    .B(_149_),
    .Y(_150_));
 sky130_fd_sc_hd__a21oi_1 _456_ (.A1(net3),
    .A2(net23),
    .B1(net55),
    .Y(_151_));
 sky130_fd_sc_hd__o22a_1 _457_ (.A1(net3),
    .A2(net23),
    .B1(_057_),
    .B2(_151_),
    .X(_152_));
 sky130_fd_sc_hd__a31o_1 _458_ (.A1(net3),
    .A2(net23),
    .A3(net56),
    .B1(_152_),
    .X(_153_));
 sky130_fd_sc_hd__a211o_1 _459_ (.A1(_058_),
    .A2(_146_),
    .B1(_150_),
    .C1(_153_),
    .X(net40));
 sky130_fd_sc_hd__and3_1 _460_ (.A(_211_),
    .B(_214_),
    .C(_131_),
    .X(_154_));
 sky130_fd_sc_hd__o21a_1 _461_ (.A1(net3),
    .A2(net23),
    .B1(_212_),
    .X(_155_));
 sky130_fd_sc_hd__o21a_1 _462_ (.A1(_220_),
    .A2(_132_),
    .B1(_154_),
    .X(_156_));
 sky130_fd_sc_hd__a211o_1 _463_ (.A1(net3),
    .A2(net23),
    .B1(_155_),
    .C1(_156_),
    .X(_157_));
 sky130_fd_sc_hd__a31o_1 _464_ (.A1(_119_),
    .A2(_133_),
    .A3(_154_),
    .B1(_157_),
    .X(_158_));
 sky130_fd_sc_hd__xnor2_1 _465_ (.A(_235_),
    .B(_158_),
    .Y(_159_));
 sky130_fd_sc_hd__o22ai_1 _466_ (.A1(_233_),
    .A2(_050_),
    .B1(net55),
    .B2(_235_),
    .Y(_160_));
 sky130_fd_sc_hd__a31o_1 _467_ (.A1(net2),
    .A2(_206_),
    .A3(_210_),
    .B1(_209_),
    .X(_161_));
 sky130_fd_sc_hd__o211a_1 _468_ (.A1(net59),
    .A2(_128_),
    .B1(_218_),
    .C1(_216_),
    .X(_162_));
 sky130_fd_sc_hd__a211o_1 _469_ (.A1(_224_),
    .A2(_032_),
    .B1(_161_),
    .C1(_162_),
    .X(_163_));
 sky130_fd_sc_hd__or2_1 _470_ (.A(_235_),
    .B(_163_),
    .X(_164_));
 sky130_fd_sc_hd__a21oi_1 _471_ (.A1(_235_),
    .A2(_163_),
    .B1(_063_),
    .Y(_165_));
 sky130_fd_sc_hd__a22o_1 _472_ (.A1(_058_),
    .A2(_159_),
    .B1(_164_),
    .B2(_165_),
    .X(_166_));
 sky130_fd_sc_hd__a211o_1 _473_ (.A1(_234_),
    .A2(_057_),
    .B1(_160_),
    .C1(_166_),
    .X(net41));
 sky130_fd_sc_hd__a21boi_2 _474_ (.A1(_234_),
    .A2(_158_),
    .B1_N(_233_),
    .Y(_167_));
 sky130_fd_sc_hd__nor2_1 _475_ (.A(_232_),
    .B(_167_),
    .Y(_168_));
 sky130_fd_sc_hd__a21o_1 _476_ (.A1(_232_),
    .A2(_167_),
    .B1(_059_),
    .X(_169_));
 sky130_fd_sc_hd__and2b_1 _477_ (.A_N(net24),
    .B(net4),
    .X(_170_));
 sky130_fd_sc_hd__a21oi_1 _478_ (.A1(_235_),
    .A2(_163_),
    .B1(_170_),
    .Y(_171_));
 sky130_fd_sc_hd__xor2_1 _479_ (.A(_232_),
    .B(_171_),
    .X(_172_));
 sky130_fd_sc_hd__and2_1 _480_ (.A(net5),
    .B(net25),
    .X(_173_));
 sky130_fd_sc_hd__nand2_1 _481_ (.A(net5),
    .B(net25),
    .Y(_174_));
 sky130_fd_sc_hd__nor2_1 _482_ (.A(net17),
    .B(_173_),
    .Y(_175_));
 sky130_fd_sc_hd__nor2_1 _483_ (.A(net5),
    .B(net25),
    .Y(_176_));
 sky130_fd_sc_hd__o22a_1 _484_ (.A1(_053_),
    .A2(_173_),
    .B1(_175_),
    .B2(_050_),
    .X(_177_));
 sky130_fd_sc_hd__o22a_1 _485_ (.A1(_063_),
    .A2(_172_),
    .B1(_176_),
    .B2(_177_),
    .X(_178_));
 sky130_fd_sc_hd__o21ai_1 _486_ (.A1(_168_),
    .A2(_169_),
    .B1(_178_),
    .Y(net42));
 sky130_fd_sc_hd__nor2_1 _487_ (.A(_167_),
    .B(_176_),
    .Y(_179_));
 sky130_fd_sc_hd__a211o_1 _488_ (.A1(_167_),
    .A2(_174_),
    .B1(_176_),
    .C1(_239_),
    .X(_180_));
 sky130_fd_sc_hd__o311a_1 _489_ (.A1(_240_),
    .A2(_173_),
    .A3(_179_),
    .B1(_180_),
    .C1(_058_),
    .X(_181_));
 sky130_fd_sc_hd__a21o_1 _490_ (.A1(_230_),
    .A2(_171_),
    .B1(_231_),
    .X(_182_));
 sky130_fd_sc_hd__xnor2_1 _491_ (.A(_239_),
    .B(_182_),
    .Y(_183_));
 sky130_fd_sc_hd__nand2_1 _492_ (.A(_238_),
    .B(_049_),
    .Y(_184_));
 sky130_fd_sc_hd__a21oi_1 _493_ (.A1(_208_),
    .A2(_237_),
    .B1(_184_),
    .Y(_185_));
 sky130_fd_sc_hd__nor2_1 _494_ (.A(_239_),
    .B(net55),
    .Y(_186_));
 sky130_fd_sc_hd__a211o_1 _495_ (.A1(_062_),
    .A2(_183_),
    .B1(_185_),
    .C1(_186_),
    .X(_187_));
 sky130_fd_sc_hd__or2_1 _496_ (.A(_181_),
    .B(_187_),
    .X(net43));
 sky130_fd_sc_hd__nand2_1 _497_ (.A(_237_),
    .B(_180_),
    .Y(_188_));
 sky130_fd_sc_hd__a21oi_1 _498_ (.A1(_237_),
    .A2(_180_),
    .B1(_228_),
    .Y(_189_));
 sky130_fd_sc_hd__a31o_1 _499_ (.A1(_228_),
    .A2(_237_),
    .A3(_180_),
    .B1(_059_),
    .X(_190_));
 sky130_fd_sc_hd__o21a_1 _500_ (.A1(_240_),
    .A2(_182_),
    .B1(_236_),
    .X(_191_));
 sky130_fd_sc_hd__or3_1 _501_ (.A(_228_),
    .B(_063_),
    .C(_191_),
    .X(_192_));
 sky130_fd_sc_hd__nor2_1 _502_ (.A(_225_),
    .B(_050_),
    .Y(_193_));
 sky130_fd_sc_hd__a221o_1 _503_ (.A1(_227_),
    .A2(_052_),
    .B1(_057_),
    .B2(_226_),
    .C1(_193_),
    .X(_194_));
 sky130_fd_sc_hd__a31oi_1 _504_ (.A1(_228_),
    .A2(_062_),
    .A3(_191_),
    .B1(_194_),
    .Y(_195_));
 sky130_fd_sc_hd__o211ai_1 _505_ (.A1(_189_),
    .A2(_190_),
    .B1(_192_),
    .C1(_195_),
    .Y(net44));
 sky130_fd_sc_hd__or4_4 _506_ (.A(net45),
    .B(net46),
    .C(net47),
    .D(net48),
    .X(_196_));
 sky130_fd_sc_hd__or4_4 _507_ (.A(net49),
    .B(net50),
    .C(net52),
    .D(_196_),
    .X(_197_));
 sky130_fd_sc_hd__or3_4 _508_ (.A(_197_),
    .B(net53),
    .C(net38),
    .X(_198_));
 sky130_fd_sc_hd__nor4_4 _509_ (.A(net51),
    .B(net39),
    .C(_198_),
    .D(net41),
    .Y(_199_));
 sky130_fd_sc_hd__nor2_1 _510_ (.A(net40),
    .B(net42),
    .Y(_200_));
 sky130_fd_sc_hd__and4bb_1 _511_ (.A_N(net43),
    .B_N(net44),
    .C(_200_),
    .D(_199_),
    .X(net54));
 sky130_fd_sc_hd__xnor2_1 _512_ (.A(net7),
    .B(_191_),
    .Y(_201_));
 sky130_fd_sc_hd__a31o_1 _513_ (.A1(_225_),
    .A2(_237_),
    .A3(_180_),
    .B1(_059_),
    .X(_202_));
 sky130_fd_sc_hd__a21oi_1 _514_ (.A1(_226_),
    .A2(_188_),
    .B1(_202_),
    .Y(_203_));
 sky130_fd_sc_hd__a31o_1 _515_ (.A1(_227_),
    .A2(_062_),
    .A3(_201_),
    .B1(_203_),
    .X(net37));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_145 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(a[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(a[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(a[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(a[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(a[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(a[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(a[1]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(a[2]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(a[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(a[4]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(a[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(a[6]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(a[7]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(a[8]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(a[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(alu_control[0]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(alu_control[1]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(alu_control[2]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(alu_control[3]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(b[0]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(b[10]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(b[11]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(b[12]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(b[13]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(b[14]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(b[15]),
    .X(net27));
 sky130_fd_sc_hd__buf_6 input28 (.A(b[1]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(b[2]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(b[3]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(b[4]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input32 (.A(b[5]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(b[6]),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(b[7]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(b[8]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(b[9]),
    .X(net36));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(overflow));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(result[0]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(result[10]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(result[11]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(result[12]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(result[13]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(result[14]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(result[15]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(result[1]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(result[2]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(result[3]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(result[4]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(result[5]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(result[6]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(result[7]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(result[8]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(result[9]));
 sky130_fd_sc_hd__buf_6 output54 (.A(net54),
    .X(zero));
 sky130_fd_sc_hd__clkbuf_4 fanout55 (.A(_053_),
    .X(net55));
 sky130_fd_sc_hd__buf_2 max_cap56 (.A(_049_),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(_214_),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(_083_),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(_217_),
    .X(net59));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_189 ();
endmodule
